module controladorVGA (CLK, R, G, B, horiz_sync, vert_sync);
	input logic CLK;
	input logic R, G, B;
	input logic horiz_sync, vert_sync;
	
	
endmodule 